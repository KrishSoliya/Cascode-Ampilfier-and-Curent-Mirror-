magic
tech scmos
timestamp 1731232218
<< nwell >>
rect -37 -22 64 63
<< ntransistor >>
rect -13 -65 -11 -55
rect 38 -65 40 -55
<< ptransistor >>
rect -13 -15 -11 33
rect 37 -15 39 33
<< ndiffusion >>
rect -20 -60 -13 -55
rect -21 -61 -13 -60
rect -21 -65 -20 -61
rect -16 -65 -13 -61
rect -11 -56 -3 -55
rect -11 -60 -8 -56
rect -4 -60 -3 -56
rect 30 -56 38 -55
rect 34 -60 38 -56
rect -11 -65 -4 -60
rect 31 -65 38 -60
rect 40 -59 42 -55
rect 46 -59 48 -55
rect 40 -60 48 -59
rect 40 -65 47 -60
<< pdiffusion >>
rect -16 29 -13 33
rect -20 -15 -13 29
rect -11 29 -8 33
rect -11 -15 -4 29
rect 34 29 37 33
rect 30 -15 37 29
rect 39 -11 46 33
rect 39 -15 42 -11
<< ndcontact >>
rect -20 -65 -16 -61
rect -8 -60 -4 -56
rect 30 -60 34 -56
rect 42 -59 46 -55
<< pdcontact >>
rect -20 29 -16 33
rect -8 29 -4 33
rect 30 29 34 33
rect 42 -15 46 -11
<< psubstratepcontact >>
rect -21 -102 -17 -98
rect 1 -103 5 -99
rect 25 -103 29 -99
rect 45 -103 49 -99
<< nsubstratencontact >>
rect -21 55 -17 59
rect -3 55 1 59
rect 20 55 24 59
rect 39 55 43 59
<< polysilicon >>
rect -13 33 -11 43
rect 37 33 39 43
rect -13 -21 -11 -15
rect 37 -22 39 -15
rect -13 -55 -11 -44
rect 38 -55 40 -44
rect -13 -73 -11 -65
rect 38 -73 40 -65
<< polycontact >>
rect -13 43 -9 47
rect 37 43 41 47
rect -13 -77 -9 -73
rect 38 -77 42 -73
<< metal1 >>
rect -36 59 61 61
rect -36 55 -21 59
rect -17 55 -3 59
rect 1 55 20 59
rect 24 55 39 59
rect 43 55 61 59
rect -36 53 61 55
rect -20 33 -16 53
rect -9 43 0 47
rect 41 43 50 47
rect -9 29 -8 33
rect -4 29 30 33
rect 46 -15 47 -11
rect 42 -55 47 -15
rect -8 -56 35 -55
rect -4 -60 30 -56
rect 34 -60 35 -56
rect 46 -58 47 -55
rect -21 -61 -16 -60
rect -21 -65 -20 -61
rect -21 -98 -16 -65
rect -9 -77 0 -73
rect 42 -77 51 -73
rect -36 -102 -21 -98
rect -17 -99 61 -98
rect -17 -102 1 -99
rect -36 -103 1 -102
rect 5 -103 25 -99
rect 29 -103 45 -99
rect 49 -103 61 -99
rect -36 -106 61 -103
<< labels >>
flabel metal1 8 54 12 58 0 FreeSans 18 0 0 0 Vdd
flabel nwell -3 43 1 47 0 FreeSans 18 0 0 0 Vbias1
flabel metal1 46 43 50 47 0 FreeSans 18 0 0 0 Vbias2
flabel metal1 -4 -77 0 -73 0 FreeSans 18 0 0 0 Vin
flabel metal1 47 -77 51 -73 0 FreeSans 18 0 0 0 Vbias3
flabel metal1 14 -103 18 -99 0 FreeSans 18 0 0 0 GND
<< end >>
